
//module shiftreg #(parameter SHIFT = 0, DATA=32)
//   (input         clk,reset,
//    input  [DATA-1:0] data_in,
//    output [DATA-1:0] data_out);

//reg [DATA-1:0] shift_array [SHIFT-1:0];

//always @(posedge clk or posedge reset) begin
//    if(reset)
//        shift_array[0] <= 0;
//    else
//        shift_array[0] <= data_in;
//end

//genvar shft;

//generate
//    for(shft=0; shft < SHIFT-1; shft=shft+1) begin: DELAY_BLOCK
//        always @(posedge clk or posedge reset) begin
//            if(reset)
//                shift_array[shft+1] <= 0;
//            else
//                shift_array[shft+1] <= shift_array[shft];
//        end
//    end
//endgenerate

//assign data_out = shift_array[SHIFT-1];

//endmodule

module shiftreg #(
    parameter SHIFT = 32,  // ��λ����
    parameter DATA  = 32   // ����λ��
) (
    input              clk, reset,      // ʱ�Ӻ��첽��λ
    input  [DATA-1:0]  data_in,         // ��������
    output [DATA-1:0]  data_out         // �������
);

generate
    if (SHIFT == 0) begin
        // �ӳ�Ϊ0��ֱ���������뵽���
        assign data_out = data_in;
    end 
    else if (SHIFT == 1) begin
        // �ӳ�Ϊ1��ֻ��һ���Ĵ���
        reg [DATA-1:0] shift_reg;
        always @(posedge clk or posedge reset) begin
            if (reset)
                shift_reg <= 0;
            else
                shift_reg <= data_in;
        end
        assign data_out = shift_reg;
    end 
    else begin
        // �ӳٴ���1��ʹ��SRLC32Eʵ��SHIFT-1����λ���ٽ�һ���Ĵ���
        wire [DATA-1:0] srl_out;
        reg [DATA-1:0] output_reg;

        genvar i;
        for (i = 0; i < DATA; i = i + 1) begin : BIT_SHIFT
            SRLC32E #(
                .INIT(32'h00000000)  // ��ʼ��ֵ
            ) srl_inst (
                .A(SHIFT-2),         // ����SHIFT-1����λ
                .CE(1'b1),           // ʼ��ʹ��
                .CLK(clk),           // ʱ��
                .D(data_in[i]),      // ��������
                .Q(srl_out[i]),      // ��λ���
                .Q31()               // δʹ��
            );
        end

        // ����Ĵ�������SRL�����֧�ָ�λ
        always @(posedge clk or posedge reset) begin
            if (reset)
                output_reg <= 0;
            else
                output_reg <= srl_out;
        end

        assign data_out = output_reg;
    end
endgenerate

endmodule

