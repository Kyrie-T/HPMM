

// read latency is 1 cc

module BROM_PRE(input             clk,
             input      [8:0]  raddr,
             output reg [11:0] dout);
// bram
(* rom_style="block" *) reg [11:0] blockrom [511:0]; 

// premultiply k_inv
always @(posedge clk) begin
    case(raddr)
    // W
    9'd0  : dout <= 12'hc7c;
    9'd1  : dout <= 12'h53a;
    9'd2  : dout <= 12'hc04;
    9'd3  : dout <= 12'h235;
    9'd4  : dout <= 12'h5d0;
    9'd5  : dout <= 12'hb6f;
    9'd6  : dout <= 12'h2bf;
    9'd7  : dout <= 12'h8af;
    9'd8  : dout <= 12'h76d;
    9'd9  : dout <= 12'haf2;
    9'd10 : dout <= 12'h3c3;
    9'd11 : dout <= 12'h32a;
    9'd12 : dout <= 12'h906;
    9'd13 : dout <= 12'h9d5;
    9'd14 : dout <= 12'h37a;
    9'd15 : dout <= 12'h9ea;
    9'd16 : dout <= 12'h244;
    9'd17 : dout <= 12'hc9a;
    9'd18 : dout <= 12'h68f;
    9'd19 : dout <= 12'h316;
    9'd20 : dout <= 12'h3fc;
    9'd21 : dout <= 12'h354;
    9'd22 : dout <= 12'h69a;
    9'd23 : dout <= 12'h893;
    9'd24 : dout <= 12'h5f ;
    9'd25 : dout <= 12'h1d7;
    9'd26 : dout <= 12'h823;
    9'd27 : dout <= 12'h48 ;
    9'd28 : dout <= 12'h523;
    9'd29 : dout <= 12'ha69;
    9'd30 : dout <= 12'h1c1;
    9'd31 : dout <= 12'h2ea;
    9'd32 : dout <= 12'h5e7;
    9'd33 : dout <= 12'h206;
    9'd34 : dout <= 12'h79 ;
    9'd35 : dout <= 12'ha4 ;
    9'd36 : dout <= 12'h24f;
    9'd37 : dout <= 12'h151;
    9'd38 : dout <= 12'h62 ;
    9'd39 : dout <= 12'hccf;
    9'd40 : dout <= 12'h68 ;
    9'd41 : dout <= 12'h33f;
    9'd42 : dout <= 12'h7d0;
    9'd43 : dout <= 12'h424;
    9'd44 : dout <= 12'h6fe;
    9'd45 : dout <= 12'h69b;
    9'd46 : dout <= 12'h36d;
    9'd47 : dout <= 12'h44e;
    9'd48 : dout <= 12'h492;
    9'd49 : dout <= 12'hc2 ;
    9'd50 : dout <= 12'h9de;
    9'd51 : dout <= 12'h792;
    9'd52 : dout <= 12'h724;
    9'd53 : dout <= 12'hc8b;
    9'd54 : dout <= 12'h948;
    9'd55 : dout <= 12'h735;
    9'd56 : dout <= 12'h337;
    9'd57 : dout <= 12'hb8f;
    9'd58 : dout <= 12'hacf;
    9'd59 : dout <= 12'h342;
    9'd60 : dout <= 12'h211;
    9'd61 : dout <= 12'h4a2;
    9'd62 : dout <= 12'hcbb;
    9'd63 : dout <= 12'h3ff;
    9'd64 : dout <= 12'h42c;
    9'd65 : dout <= 12'had4;
    9'd66 : dout <= 12'h935;
    9'd67 : dout <= 12'hb83;
    9'd68 : dout <= 12'h7c9;
    9'd69 : dout <= 12'hc51;
    9'd70 : dout <= 12'h7ac;
    9'd71 : dout <= 12'h494;
    9'd72 : dout <= 12'h934;
    9'd73 : dout <= 12'h404;
    9'd74 : dout <= 12'hbef;
    9'd75 : dout <= 12'h1c6;
    9'd76 : dout <= 12'ha5b;
    9'd77 : dout <= 12'hb19;
    9'd78 : dout <= 12'h716;
    9'd79 : dout <= 12'hc7e;
    9'd80 : dout <= 12'hc82;
    9'd81 : dout <= 12'h62a;
    9'd82 : dout <= 12'h777;
    9'd83 : dout <= 12'h72 ;
    9'd84 : dout <= 12'h2b7;
    9'd85 : dout <= 12'h490;
    9'd86 : dout <= 12'h832;
    9'd87 : dout <= 12'h2b8;
    9'd88 : dout <= 12'h64f;
    9'd89 : dout <= 12'h545;
    9'd90 : dout <= 12'h849;
    9'd91 : dout <= 12'h4c8;
    9'd92 : dout <= 12'h94d;
    9'd93 : dout <= 12'h7ec;
    9'd94 : dout <= 12'h3cf;
    9'd95 : dout <= 12'ha87;
    9'd96 : dout <= 12'h950;
    9'd97 : dout <= 12'h864;
    9'd98 : dout <= 12'h809;
    9'd99 : dout <= 12'hae4;
    9'd100: dout <= 12'h3c ;
    9'd101: dout <= 12'h960;
    9'd102: dout <= 12'h682;
    9'd103: dout <= 12'h9af;
    9'd104: dout <= 12'h6e8;
    9'd105: dout <= 12'h32b;
    9'd106: dout <= 12'h2c6;
    9'd107: dout <= 12'h55f;
    9'd108: dout <= 12'h1d5;
    9'd109: dout <= 12'h843;
    9'd110: dout <= 12'h639;
    9'd111: dout <= 12'h829;
    9'd112: dout <= 12'hcad;
    9'd113: dout <= 12'hce2;
    9'd114: dout <= 12'hbb2;
    9'd115: dout <= 12'hba9;
    9'd116: dout <= 12'h45b;
    9'd117: dout <= 12'h52b;
    9'd118: dout <= 12'h1bc;
    9'd119: dout <= 12'h57c;
    9'd120: dout <= 12'h2a3;
    9'd121: dout <= 12'h170;
    9'd122: dout <= 12'h1b1;
    9'd123: dout <= 12'h35e;
    9'd124: dout <= 12'h91f;
    9'd125: dout <= 12'hbc ;
    9'd126: dout <= 12'h85b;
    
    // WINV
    9'd127: dout <= 12'h4a6;
    9'd128: dout <= 12'hc45;
    9'd129: dout <= 12'h3e2;
    9'd130: dout <= 12'h9a3;
    9'd131: dout <= 12'hb50;
    9'd132: dout <= 12'hb91;
    9'd133: dout <= 12'ha5e;
    9'd134: dout <= 12'h785;
    9'd135: dout <= 12'hb45;
    9'd136: dout <= 12'h7d6;
    9'd137: dout <= 12'h8a6;
    9'd138: dout <= 12'h158;
    9'd139: dout <= 12'h14f;
    9'd140: dout <= 12'h1f ;
    9'd141: dout <= 12'h54 ;
    9'd142: dout <= 12'h4d8;
    9'd143: dout <= 12'h6c8;
    9'd144: dout <= 12'h4be;
    9'd145: dout <= 12'hb2c;
    9'd146: dout <= 12'h7a2;
    9'd147: dout <= 12'ha3b;
    9'd148: dout <= 12'h9d6;
    9'd149: dout <= 12'h619;
    9'd150: dout <= 12'h352;
    9'd151: dout <= 12'h67f;
    9'd152: dout <= 12'h3a1;
    9'd153: dout <= 12'hcc5;
    9'd154: dout <= 12'h21d;
    9'd155: dout <= 12'h4f8;
    9'd156: dout <= 12'h49d;
    9'd157: dout <= 12'h3b1;
    9'd158: dout <= 12'h27a;
    9'd159: dout <= 12'h932;
    9'd160: dout <= 12'h515;
    9'd161: dout <= 12'h3b4;
    9'd162: dout <= 12'h839;
    9'd163: dout <= 12'h4b8;
    9'd164: dout <= 12'h7bc;
    9'd165: dout <= 12'h6b2;
    9'd166: dout <= 12'ha49;
    9'd167: dout <= 12'h4cf;
    9'd168: dout <= 12'h871;
    9'd169: dout <= 12'ha4a;
    9'd170: dout <= 12'hc8f;
    9'd171: dout <= 12'h58a;
    9'd172: dout <= 12'h6d7;
    9'd173: dout <= 12'h7f ;
    9'd174: dout <= 12'h83 ;
    9'd175: dout <= 12'h5eb;
    9'd176: dout <= 12'h1e8;
    9'd177: dout <= 12'h2a6;
    9'd178: dout <= 12'hb3b;
    9'd179: dout <= 12'h112;
    9'd180: dout <= 12'h8fd;
    9'd181: dout <= 12'h3cd;
    9'd182: dout <= 12'h86d;
    9'd183: dout <= 12'h555;
    9'd184: dout <= 12'hb0 ;
    9'd185: dout <= 12'h538;
    9'd186: dout <= 12'h17e;
    9'd187: dout <= 12'h3cc;
    9'd188: dout <= 12'h22d;
    9'd189: dout <= 12'h8d5;
    9'd190: dout <= 12'h902;
    9'd191: dout <= 12'h46 ;
    9'd192: dout <= 12'h85f;
    9'd193: dout <= 12'haf0;
    9'd194: dout <= 12'h9bf;
    9'd195: dout <= 12'h232;
    9'd196: dout <= 12'h172;
    9'd197: dout <= 12'h9ca;
    9'd198: dout <= 12'h5cc;
    9'd199: dout <= 12'h3b9;
    9'd200: dout <= 12'h76 ;
    9'd201: dout <= 12'h5dd;
    9'd202: dout <= 12'h56f;
    9'd203: dout <= 12'h323;
    9'd204: dout <= 12'hc3f;
    9'd205: dout <= 12'h86f;
    9'd206: dout <= 12'h8b3;
    9'd207: dout <= 12'h994;
    9'd208: dout <= 12'h666;
    9'd209: dout <= 12'h603;
    9'd210: dout <= 12'h8dd;
    9'd211: dout <= 12'h531;
    9'd212: dout <= 12'h9c2;
    9'd213: dout <= 12'hc99;
    9'd214: dout <= 12'h32 ;
    9'd215: dout <= 12'hc9f;
    9'd216: dout <= 12'hbb0;
    9'd217: dout <= 12'hab2;
    9'd218: dout <= 12'hc5d;
    9'd219: dout <= 12'hc88;
    9'd220: dout <= 12'hafb;
    9'd221: dout <= 12'h71a;
    9'd222: dout <= 12'ha17;
    9'd223: dout <= 12'hb40;
    9'd224: dout <= 12'h298;
    9'd225: dout <= 12'h7de;
    9'd226: dout <= 12'hcb9;
    9'd227: dout <= 12'h4de;
    9'd228: dout <= 12'hb2a;
    9'd229: dout <= 12'hca2;
    9'd230: dout <= 12'h46e;
    9'd231: dout <= 12'h667;
    9'd232: dout <= 12'h9ad;
    9'd233: dout <= 12'h905;
    9'd234: dout <= 12'h9eb;
    9'd235: dout <= 12'h672;
    9'd236: dout <= 12'h67 ;
    9'd237: dout <= 12'habd;
    9'd238: dout <= 12'h317;
    9'd239: dout <= 12'h987;
    9'd240: dout <= 12'h32c;
    9'd241: dout <= 12'h3fb;
    9'd242: dout <= 12'h9d7;
    9'd243: dout <= 12'h93e;
    9'd244: dout <= 12'h20f;
    9'd245: dout <= 12'h594;
    9'd246: dout <= 12'h452;
    9'd247: dout <= 12'ha42;
    9'd248: dout <= 12'h192;
    9'd249: dout <= 12'h731;
    9'd250: dout <= 12'hacc;
    9'd251: dout <= 12'hfd ;
    9'd252: dout <= 12'h7c7;
    9'd253: dout <= 12'h85 ;
    // W MULT
    9'd254: dout <= 12'h3ff;
    9'd255: dout <= 12'h902;
    9'd256: dout <= 12'h42c;
    9'd257: dout <= 12'h8d5;
    9'd258: dout <= 12'had4;
    9'd259: dout <= 12'h22d;
    9'd260: dout <= 12'h935;
    9'd261: dout <= 12'h3cc;
    9'd262: dout <= 12'hb83;
    9'd263: dout <= 12'h17e;
    9'd264: dout <= 12'h7c9;
    9'd265: dout <= 12'h538;
    9'd266: dout <= 12'hc51;
    9'd267: dout <= 12'hb0 ;
    9'd268: dout <= 12'h7ac;
    9'd269: dout <= 12'h555;
    9'd270: dout <= 12'h494;
    9'd271: dout <= 12'h86d;
    9'd272: dout <= 12'h934;
    9'd273: dout <= 12'h3cd;
    9'd274: dout <= 12'h404;
    9'd275: dout <= 12'h8fd;
    9'd276: dout <= 12'hbef;
    9'd277: dout <= 12'h112;
    9'd278: dout <= 12'h1c6;
    9'd279: dout <= 12'hb3b;
    9'd280: dout <= 12'ha5b;
    9'd281: dout <= 12'h2a6;
    9'd282: dout <= 12'hb19;
    9'd283: dout <= 12'h1e8;
    9'd284: dout <= 12'h716;
    9'd285: dout <= 12'h5eb;
    9'd286: dout <= 12'hc7e;
    9'd287: dout <= 12'h83 ;
    9'd288: dout <= 12'hc82;
    9'd289: dout <= 12'h7f ;
    9'd290: dout <= 12'h62a;
    9'd291: dout <= 12'h6d7;
    9'd292: dout <= 12'h777;
    9'd293: dout <= 12'h58a;
    9'd294: dout <= 12'h72 ;
    9'd295: dout <= 12'hc8f;
    9'd296: dout <= 12'h2b7;
    9'd297: dout <= 12'ha4a;
    9'd298: dout <= 12'h490;
    9'd299: dout <= 12'h871;
    9'd300: dout <= 12'h832;
    9'd301: dout <= 12'h4cf;
    9'd302: dout <= 12'h2b8;
    9'd303: dout <= 12'ha49;
    9'd304: dout <= 12'h64f;
    9'd305: dout <= 12'h6b2;
    9'd306: dout <= 12'h545;
    9'd307: dout <= 12'h7bc;
    9'd308: dout <= 12'h849;
    9'd309: dout <= 12'h4b8;
    9'd310: dout <= 12'h4c8;
    9'd311: dout <= 12'h839;
    9'd312: dout <= 12'h94d;
    9'd313: dout <= 12'h3b4;
    9'd314: dout <= 12'h7ec;
    9'd315: dout <= 12'h515;
    9'd316: dout <= 12'h3cf;
    9'd317: dout <= 12'h932;
    9'd318: dout <= 12'ha87;
    9'd319: dout <= 12'h27a;
    9'd320: dout <= 12'h950;
    9'd321: dout <= 12'h3b1;
    9'd322: dout <= 12'h864;
    9'd323: dout <= 12'h49d;
    9'd324: dout <= 12'h809;
    9'd325: dout <= 12'h4f8;
    9'd326: dout <= 12'hae4;
    9'd327: dout <= 12'h21d;
    9'd328: dout <= 12'h3c ;
    9'd329: dout <= 12'hcc5;
    9'd330: dout <= 12'h960;
    9'd331: dout <= 12'h3a1;
    9'd332: dout <= 12'h682;
    9'd333: dout <= 12'h67f;
    9'd334: dout <= 12'h9af;
    9'd335: dout <= 12'h352;
    9'd336: dout <= 12'h6e8;
    9'd337: dout <= 12'h619;
    9'd338: dout <= 12'h32b;
    9'd339: dout <= 12'h9d6;
    9'd340: dout <= 12'h2c6;
    9'd341: dout <= 12'ha3b;
    9'd342: dout <= 12'h55f;
    9'd343: dout <= 12'h7a2;
    9'd344: dout <= 12'h1d5;
    9'd345: dout <= 12'hb2c;
    9'd346: dout <= 12'h843;
    9'd347: dout <= 12'h4be;
    9'd348: dout <= 12'h639;
    9'd349: dout <= 12'h6c8;
    9'd350: dout <= 12'h829;
    9'd351: dout <= 12'h4d8;
    9'd352: dout <= 12'hcad;
    9'd353: dout <= 12'h54 ;
    9'd354: dout <= 12'hce2;
    9'd355: dout <= 12'h1f ;
    9'd356: dout <= 12'hbb2;
    9'd357: dout <= 12'h14f;
    9'd358: dout <= 12'hba9;
    9'd359: dout <= 12'h158;
    9'd360: dout <= 12'h45b;
    9'd361: dout <= 12'h8a6;
    9'd362: dout <= 12'h52b;
    9'd363: dout <= 12'h7d6;
    9'd364: dout <= 12'h1bc;
    9'd365: dout <= 12'hb45;
    9'd366: dout <= 12'h57c;
    9'd367: dout <= 12'h785;
    9'd368: dout <= 12'h2a3;
    9'd369: dout <= 12'ha5e;
    9'd370: dout <= 12'h170;
    9'd371: dout <= 12'hb91;
    9'd372: dout <= 12'h1b1;
    9'd373: dout <= 12'hb50;
    9'd374: dout <= 12'h35e;
    9'd375: dout <= 12'h9a3;
    9'd376: dout <= 12'h91f;
    9'd377: dout <= 12'h3e2;
    9'd378: dout <= 12'hbc ;
    9'd379: dout <= 12'hc45;
    9'd380: dout <= 12'h85b;
    9'd381: dout <= 12'h4a6;
    default: dout <= 12'h0;
    endcase
end

endmodule
