
//module modsub(input [11:0] A,B,
//              output reg [11:0] C);

//reg signed [12:0] R;
//reg signed [12:0] Rq;

//always @(*) begin
//    R = A - B;
//    if (R[12] == 0) begin // R >= 0
//        C = R[11:0];
//    end else begin // R < 0
//        Rq= R + 13'd3329;
//        C = Rq[11:0];
//    end
//end

//endmodule

module modsub #(
    parameter LOGQ       = 12,            // ����λ��Ϊ 12 λ
    parameter [LOGQ:0] Q_VALUE = 13'd3329 // �̶�ģ��Ϊ 3329
) (
    input  [LOGQ-1:0] a,   // ���� a��12 λ��
    input  [LOGQ-1:0] b,   // ���� b��12 λ��
    output [LOGQ-1:0] c    // ��� c��12 λ��
);

// ------------------------------------------
// ����߼�ʵ�֣���ʱ�ӺͼĴ�����
// ------------------------------------------
wire signed [LOGQ:0]   msub;      // ��ʱ���������13 λ�з�������
wire signed [LOGQ:0] msub_q; // ����ģ������з��Ž����13 λ�з�������

assign msub = a + ~b + 1;                // ���� a - b��13 λ�з�������
assign msub_q = msub + Q_VALUE;     // ����ģ�� 3329��13 λ�з�������

// ���ѡ���� msub �Ǹ���ȡ����������������ģ�����
assign c = (msub[LOGQ] == 0) ? msub[LOGQ-1:0] : msub_q[LOGQ-1:0];

endmodule

//module modsub #(
//    parameter LOGQ       = 12,            // ����λ��Ϊ 12 λ
//    parameter [LOGQ:0] Q_VALUE = 13'd3329 // �̶�ģ��Ϊ 3329
//) (
//    input  [LOGQ-1:0] a,   // ���� a��12 λ��
//    input  [LOGQ-1:0] b,   // ���� b��12 λ��
//    output [LOGQ-1:0] c    // ��� c��12 λ��
//);

//wire signed [LOGQ:0] msub = a - b;       // ��һ������13 λ�з�������
//wire signed [LOGQ:0] sub_result = (msub < 0) ? msub + Q_VALUE : msub;
//assign c = sub_result[LOGQ-1:0];         // ȡ�� 12 λ

//endmodule
