
// module modadd(input [11:0] A,B,
//               output[11:0] C);

// wire        [12:0] R;
// wire signed [13:0] Rq;

// assign R = A + B;
// assign Rq= R - 13'd3329;

// assign C = (Rq[13] == 0) ? Rq[11:0] : R[11:0];

// endmodule

module modadd #(
    parameter LOGQ       = 12,            // ����λ��Ϊ 12 λ����Ӧ 12 λ���������
    parameter [LOGQ:0] Q_VALUE = 13'd3329 // �̶�ģ��Ϊ 3329���� 13 λ�洢��
) (
    input  [LOGQ-1:0] a,   // ���� a��12 λ��
    input  [LOGQ-1:0] b,   // ���� b��12 λ��
    output [LOGQ-1:0] c    // ��� c��12 λ��
);

// ------------------------------------------
// ����߼�ʵ�֣���ʱ�ӺͼĴ�����
// ------------------------------------------
wire [LOGQ:0]   madd;      // ��ʱ�ӷ������13 λ��
wire signed [LOGQ+1:0] madd_q; // ģ������з��Ž����14 λ��

assign madd = a + b;                // ���� a + b��13 λ��
assign madd_q = madd - Q_VALUE;     // ��ȥģ�� 3329��14 λ�з�������

// ���ѡ���� madd_q �Ǹ���ȡ�� 12 λ���������ӷ����
assign c = (madd_q[LOGQ+1] == 0) ? madd_q[LOGQ-1:0] : madd[LOGQ-1:0];

endmodule

//module modadd #(
//    parameter LOGQ       = 12,
//    parameter [LOGQ:0] Q_VALUE = 13'd3329
//) (
//    input  [LOGQ-1:0] a,
//    input  [LOGQ-1:0] b,
//    output [LOGQ-1:0] c
//);

//wire [LOGQ:0] madd = a + b;            // ��һ�ӷ�
//wire [LOGQ:0] sub_result = (madd >= Q_VALUE) ? madd - Q_VALUE : madd;
//assign c = sub_result[LOGQ-1:0];       // ȡ�� 12 λ

//endmodule
